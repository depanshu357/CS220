module full_sub(a,b,cin,cout,crr);
    input a,b,cin;
    output cout,crr;
    
    and and1(crr,cin,~a);
    and and1()
    
    
endmodule